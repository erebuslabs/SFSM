module fsm_rd_094_s (RST, CLK, ptext, rtext);
//user interface
	input RST, CLK;
	input [1:0] ptext;
	output[2:0] rtext;
	reg [2:0] rtext;
//STATE ASSIGNMENTS
	`include "fsm_rd_094_s_stassign.v";
   //process modeling state register
   always @ (posedge RST or posedge CLK) begin
      if( RST == 1) begin
	 State <= st1;
	 //NextState <= WT;
      end
      else
	State <= NextState;
   end
   always @ (State or ptext) begin
      case ( State )
	  st1: begin
		if(1)
 		  NextState <= st2;
		rtext <= 'b000;
	  end
	  st2: begin
		if(ptext[1] == 1 )
 		  NextState <= st3;
		else if(ptext[1] == 0 )
 		  NextState <= st2_n;
		rtext <= 'b000;
	  end
	  st2_n: begin
		if(ptext[1] == 1 )
 		  NextState <= st3;
		else if(ptext[1] == 0 )
 		  NextState <= st2;
		rtext <= 'b000;
	  end
	  st3: begin
		if(1)
 		  NextState <= st4;
		rtext <= 'b010;
	  end
	  st4: begin
		if(1)
 		  NextState <= st5;
		rtext <= 'b000;
	  end
	  st5: begin
		if(1)
 		  NextState <= st6;
		rtext <= 'b000;
	  end
	  st6: begin
		if(1)
 		  NextState <= st7;
		rtext <= 'b100;
	  end
	  st7: begin
		if(1)
 		  NextState <= st1;
		rtext <= 'b100;
	  end
      endcase // case ( State )
   end // always @ (State or ptext)   
endmodule // fsm
